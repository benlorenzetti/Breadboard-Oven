*** heat-model.cir ***
; Nodes:
; gnd, atm, bulkAir, interiorFrame, exteriorFrame, elementSurface, hotBolts, boltRadiators
;
; Nichrome Wire Heating Element Parameters:
.param Diameter=32	; [0.001 in]
.param Length=240	; [in]
.param Relement={(Length/12)*675/(Diameter*Diameter)}	; [Ohms]
.param wattage={(120*120)/Relement}
.param Volume={3.1415*Diameter*Diameter*0.000001*0.25*Length}	; [in^3]
.param SurfaceArea={3.1415*0.001*Diameter*Length*0.0254*0.0254}	; [m^2]
.param Cnichrome={0.1251*450*Volume}	; [J/K]
.param Rnichrome={0.1/SurfaceArea}	; [K/W]
;
; Frame Parameters:
.param chamberVolume=360
.param Rinsulation=3.8
.param frameWidth=4.76mm
.param Rxframe=0.0181
.param Cxframe=798.3k
.param RexteriorFrame=6.06

.param hangLength=50mm

Vroomtemp atm gnd DC 20

*Ielement atm elementSurface PULSE(0 {wattage} 1s 1ns 1ns 100s 100s)
* (initial_value, pulsed_value, delay_time, rise_time, fall_time, pulse_width, period)
Velement elementSurface atm PULSE(0 800 1s 1ns 1ns 100s 100s)

Celement elementSurface atm {Cnichrome}
RnichromeSuface elementSurface bulkAir {Rnichrome}

Rinsulate bulkAir interiorFrame {Rinsulation}

Ualuminumframe interiorFrame exteriorFrame gnd frameModel L={frameWidth}
.MODEL frameModel URC RPERL={Rxframe} CPERL={Cxframe}

Rframe exteriorFrame atm {RexteriorFrame}

Xairheatcapacity bulkAir atm varCap VOLUME={chamberVolume}

.subckt varCap n1 n2 VOLUME=360 ; inches squared
B1 n1 int2 V=273.16*(exp((v(int))/(5.8413*{VOLUME}))-1)
Vammeter int2 n2 0
F1 gnd int Vammeter 1
C1 int gnd 1
.ends varCap

.control
tran 10ms 100s; tstep, tstop
plot v(elementSurface) v(bulkAir) ;v(interiorFrame) v(exteriorFrame)

.end
